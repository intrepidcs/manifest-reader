library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package empty_pkg is

end package empty_pkg;

package body empty_pkg is

end package body empty_pkg;
